`timescale 1ns / 1ps

module datapath_debug_tb;

    // Inputs
    reg clk;
    reg rst_n;

    // Outputs
    wire [31:0] aluResult;
    wire [1:0] alu_op;
    wire [31:0] instr;
    wire [31:0] signImm;
	 wire jump;
	 wire ifbranch;

    // Instantiate the Unit Under Test (UUT)
    datapath_debug uut (
        .clk(clk),
        .rst_n(rst_n),
        .aluResult(aluResult),
        .alu_op(alu_op),
        .instr(instr),
        .signImm(signImm),
		  .jump(jump),
		  .ifbranch(ifbranch)
    );

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 100 MHz clock (10 ns period)
    end

    // Stimulus process
    initial begin
        // Initialize Inputs
        rst_n = 0;

        // Apply reset
        #20;
        rst_n = 1;

        // Run simulation for 200 cycles to observe behavior
        #2000;

        // Stop simulation
        $display("Simulation finished at time %0t", $time);
        $finish;
    end

    // Monitor outputs
    initial begin
        $monitor("Time=%0t, rst_n=%b, instr=%h, aluResult=%d, alu_op=%b, signImm=%d,  jump=%b,  ifbranch=%b",
                 $time, rst_n, instr, aluResult, alu_op, signImm, jump, ifbranch);
    end

endmodule