library verilog;
use verilog.vl_types.all;
entity tb_gpio is
end tb_gpio;
