library verilog;
use verilog.vl_types.all;
entity datapath_debug_vlg_vec_tst is
end datapath_debug_vlg_vec_tst;
